library IEEE;
use IEEE.std_logic_1164.all;  
use IEEE.numeric_std.all;     

use work.pRegisterBus.all;

package pReg_mikey is

   -- range 0xFC00 .. 0xFDFF
   --   (                                  adr      upper    lower    size   default   accesstype)
   constant TIM0BKUP     : regmap_type := (16#100#,   7,      0,        1,        0,   readwrite);
   constant TIM0CTLA     : regmap_type := (16#101#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM0CNT      : regmap_type := (16#102#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM0CTLB     : regmap_type := (16#103#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM1BKUP     : regmap_type := (16#104#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM1CTLA     : regmap_type := (16#105#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM1CNT      : regmap_type := (16#106#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM1CTLB     : regmap_type := (16#107#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM2BKUP     : regmap_type := (16#108#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM2CTLA     : regmap_type := (16#109#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM2CNT      : regmap_type := (16#10a#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM2CTLB     : regmap_type := (16#10b#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM3BKUP     : regmap_type := (16#10c#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM3CTLA     : regmap_type := (16#10d#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM3CNT      : regmap_type := (16#10e#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM3CTLB     : regmap_type := (16#10f#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM4BKUP     : regmap_type := (16#110#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM4CTLA     : regmap_type := (16#111#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM4CNT      : regmap_type := (16#112#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM4CTLB     : regmap_type := (16#113#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM5BKUP     : regmap_type := (16#114#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM5CTLA     : regmap_type := (16#115#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM5CNT      : regmap_type := (16#116#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM5CTLB     : regmap_type := (16#117#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM6BKUP     : regmap_type := (16#118#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM6CTLA     : regmap_type := (16#119#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM6CNT      : regmap_type := (16#11a#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM6CTLB     : regmap_type := (16#11b#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM7BKUP     : regmap_type := (16#11c#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM7CTLA     : regmap_type := (16#11d#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM7CNT      : regmap_type := (16#11e#,   7,      0,        1,        0,   readwrite);                                              
   constant TIM7CTLB     : regmap_type := (16#11f#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD0VOL      : regmap_type := (16#120#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD0SHFTFB   : regmap_type := (16#121#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD0OUTVAL   : regmap_type := (16#122#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD0L8SHFT   : regmap_type := (16#123#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD0TBACK    : regmap_type := (16#124#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD0CTL      : regmap_type := (16#125#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD0COUNT    : regmap_type := (16#126#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD0MISC     : regmap_type := (16#127#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD1VOL      : regmap_type := (16#128#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD1SHFTFB   : regmap_type := (16#129#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD1OUTVAL   : regmap_type := (16#12a#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD1L8SHFT   : regmap_type := (16#12b#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD1TBACK    : regmap_type := (16#12c#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD1CTL      : regmap_type := (16#12d#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD1COUNT    : regmap_type := (16#12e#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD1MISC     : regmap_type := (16#12f#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD2VOL      : regmap_type := (16#130#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD2SHFTFB   : regmap_type := (16#131#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD2OUTVAL   : regmap_type := (16#132#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD2L8SHFT   : regmap_type := (16#133#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD2TBACK    : regmap_type := (16#134#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD2CTL      : regmap_type := (16#135#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD2COUNT    : regmap_type := (16#136#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD2MISC     : regmap_type := (16#137#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD3VOL      : regmap_type := (16#138#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD3SHFTFB   : regmap_type := (16#139#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD3OUTVAL   : regmap_type := (16#13a#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD3L8SHFT   : regmap_type := (16#13b#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD3TBACK    : regmap_type := (16#13c#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD3CTL      : regmap_type := (16#13d#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD3COUNT    : regmap_type := (16#13e#,   7,      0,        1,        0,   readwrite);                                              
   constant AUD3MISC     : regmap_type := (16#13f#,   7,      0,        1,        0,   readwrite);                                              
   constant ATTEN_A      : regmap_type := (16#140#,   7,      0,        1,        0,   readwrite);                                              
   constant ATTEN_B      : regmap_type := (16#141#,   7,      0,        1,        0,   readwrite);                                              
   constant ATTEN_C      : regmap_type := (16#142#,   7,      0,        1,        0,   readwrite);                                              
   constant ATTEN_D      : regmap_type := (16#143#,   7,      0,        1,        0,   readwrite);                                              
   constant MPAN         : regmap_type := (16#144#,   7,      0,        1,        0,   readwrite);                                              
   constant MSTEREO      : regmap_type := (16#150#,   7,      0,        1,        0,   readwrite);                                              
   constant INTRST       : regmap_type := (16#180#,   7,      0,        1,        0,   readwrite);                                              
   constant INTSET       : regmap_type := (16#181#,   7,      0,        1,        0,   readwrite);                                              
   constant MAGRDY0      : regmap_type := (16#184#,   7,      0,        1,        0,   readwrite);                                              
   constant MAGRDY1      : regmap_type := (16#185#,   7,      0,        1,        0,   readwrite);                                              
   constant AUDIN        : regmap_type := (16#186#,   7,      0,        1,      128,   readwrite);                                              
   constant SYSCTL1      : regmap_type := (16#187#,   7,      0,        1,        0,   readwrite);                                              
   constant MIKEYHREV    : regmap_type := (16#188#,   7,      0,        1,        0,   readwrite);                                              
   constant MIKEYSREV    : regmap_type := (16#189#,   7,      0,        1,        0,   readwrite);                                              
   constant IODIR        : regmap_type := (16#18a#,   7,      0,        1,        0,   readwrite);                                              
   constant IODAT        : regmap_type := (16#18b#,   7,      0,        1,        0,   readwrite);                                              
   constant SERCTL       : regmap_type := (16#18c#,   7,      0,        1,        0,   readwrite);                                              
   constant SERDAT       : regmap_type := (16#18d#,   7,      0,        1,        0,   readwrite);                                              
   constant SDONEACK     : regmap_type := (16#190#,   7,      0,        1,        0,   readwrite);                                              
   constant CPUSLEEP     : regmap_type := (16#191#,   7,      0,        1,        0,   readwrite);                                              
   constant DISPCTL      : regmap_type := (16#192#,   7,      0,        1,        0,   readwrite);                                              
   constant PBKUP        : regmap_type := (16#193#,   7,      0,        1,        0,   readwrite);                                              
   constant DISPADR      : regmap_type := (16#194#,   7,      0,        1,        0,   readwrite);                                              
   constant DISPADRL     : regmap_type := (16#194#,   7,      0,        1,        0,   readwrite);                                              
   constant DISPADRH     : regmap_type := (16#195#,   7,      0,        1,        0,   readwrite);                                              
   constant Mtest0       : regmap_type := (16#19c#,   7,      0,        1,        0,   readwrite);                                              
   constant Mtest1       : regmap_type := (16#19d#,   7,      0,        1,        0,   readwrite);                                              
   constant Mtest2       : regmap_type := (16#19e#,   7,      0,        1,        0,   readwrite);                                              
   constant GREEN        : regmap_type := (16#1a0#,   3,      0,       16,        0,   readwrite);                                                                       
   constant BLUERED      : regmap_type := (16#1b0#,   7,      0,       16,        0,   readwrite);                                                                                     
   constant MMAPCTL      : regmap_type := (16#1f9#,   7,      0,        1,        0,   readwrite);                                              
   constant CPUNMI       : regmap_type := (16#1fa#,   7,      0,        1,        0,   readwrite);                                              
   constant CPUNMIL      : regmap_type := (16#1fa#,   7,      0,        1,        0,   readwrite);                                              
   constant CPUNMIH      : regmap_type := (16#1fb#,   7,      0,        1,        0,   readwrite);                                              
   constant CPURESET     : regmap_type := (16#1fc#,   7,      0,        1,        0,   readwrite);                                              
   constant CPURESETL    : regmap_type := (16#1fc#,   7,      0,        1,        0,   readwrite);                                              
   constant CPURESETH    : regmap_type := (16#1fd#,   7,      0,        1,        0,   readwrite);                                              
   constant CPUINT       : regmap_type := (16#1fe#,   7,      0,        1,        0,   readwrite);                                              
   constant CPUINTL      : regmap_type := (16#1fe#,   7,      0,        1,        0,   readwrite);                                              
   constant CPUINTH      : regmap_type := (16#1ff#,   7,      0,        1,        0,   readwrite);                                              
   
end package;
